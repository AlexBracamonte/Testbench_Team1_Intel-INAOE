module Xor_Gate(a,b,q);
  input a,b;
  output q;
  
  xor(q,a,b);
endmodule